magic
tech scmos
timestamp 1636647610
<< nwell >>
rect -16 -10 39 9
<< ntransistor >>
rect -5 -35 -3 -31
rect 5 -35 7 -31
rect 26 -35 28 -31
<< ptransistor >>
rect -5 -1 -3 3
rect 5 -1 7 3
rect 26 -1 28 3
<< ndiffusion >>
rect -7 -35 -5 -31
rect -3 -35 5 -31
rect 7 -35 9 -31
rect 25 -35 26 -31
rect 28 -35 29 -31
<< pdiffusion >>
rect -6 -1 -5 3
rect -3 -1 -1 3
rect 3 -1 5 3
rect 7 -1 8 3
rect 25 -1 26 3
rect 28 -1 29 3
<< ndcontact >>
rect -11 -35 -7 -31
rect 9 -35 13 -31
rect 21 -35 25 -31
rect 29 -35 33 -31
<< pdcontact >>
rect -10 -1 -6 3
rect -1 -1 3 3
rect 8 -1 12 3
rect 21 -1 25 3
rect 29 -1 33 3
<< polysilicon >>
rect -5 3 -3 8
rect 5 3 7 8
rect 26 3 28 8
rect -5 -31 -3 -1
rect 5 -31 7 -1
rect 26 -31 28 -1
rect -5 -38 -3 -35
rect 5 -38 7 -35
rect 26 -38 28 -35
<< polycontact >>
rect -9 -19 -5 -15
rect 1 -28 5 -24
rect 22 -20 26 -16
<< metal1 >>
rect -10 12 39 16
rect -10 3 -6 12
rect 8 3 12 12
rect 21 3 25 12
rect -10 -19 -9 -15
rect -1 -16 3 -1
rect 29 -14 33 -1
rect -1 -20 22 -16
rect 29 -18 42 -14
rect 0 -28 1 -24
rect 9 -31 13 -20
rect 29 -31 33 -18
rect -11 -39 -7 -35
rect 21 -39 25 -35
rect -11 -43 39 -39
<< labels >>
rlabel metal1 42 -18 42 -14 7 F
rlabel metal1 39 12 39 16 6 VDD
rlabel metal1 39 -43 39 -39 8 GND
rlabel metal1 -10 -19 -10 -15 1 A
rlabel metal1 0 -28 0 -24 1 B
<< end >>
