magic
tech scmos
timestamp 1639079816
<< nwell >>
rect -47 6 54 16
<< polysilicon >>
rect -15 13 -11 15
rect -7 13 -3 15
rect 19 13 26 15
rect -39 11 -37 13
rect -31 11 -29 13
rect -14 11 -12 13
rect -6 11 -4 13
rect 11 11 13 13
rect 19 11 21 13
rect 40 11 42 13
rect -39 -3 -37 7
rect -31 -3 -29 7
rect -14 -3 -12 7
rect -6 -3 -4 7
rect 11 -3 13 7
rect 19 -3 21 7
rect 40 -3 42 7
rect -39 -9 -37 -7
rect -31 -9 -29 -7
rect -14 -9 -12 -7
rect -6 -9 -4 -7
rect 11 -9 13 -7
rect 19 -9 21 -7
rect 40 -9 42 -7
<< ndiffusion >>
rect -40 -7 -39 -3
rect -37 -7 -31 -3
rect -29 -7 -28 -3
rect -15 -7 -14 -3
rect -12 -7 -6 -3
rect -4 -7 -3 -3
rect 10 -7 11 -3
rect 13 -7 19 -3
rect 21 -7 22 -3
rect 35 -7 40 -3
rect 42 -7 47 -3
<< pdiffusion >>
rect -40 7 -39 11
rect -37 7 -36 11
rect -32 7 -31 11
rect -29 7 -28 11
rect -15 7 -14 11
rect -12 7 -11 11
rect -7 7 -6 11
rect -4 7 -3 11
rect 10 7 11 11
rect 13 7 14 11
rect 18 7 19 11
rect 21 7 22 11
rect 35 7 40 11
rect 42 7 47 11
<< metal1 >>
rect -36 15 -15 19
rect -3 15 18 19
rect 26 15 51 19
rect -36 11 -32 15
rect 14 11 18 15
rect 47 11 51 15
rect -36 4 -32 7
rect -11 4 -7 7
rect 14 4 18 7
rect -36 0 -24 4
rect -11 0 1 4
rect 14 0 26 4
rect -28 -3 -24 0
rect -3 -3 1 0
rect 22 -3 26 0
rect 47 -3 51 7
rect -44 -14 -41 -7
rect -19 -14 -16 -7
rect 6 -14 9 -7
rect 31 -14 34 -7
rect -44 -17 51 -14
<< ntransistor >>
rect -39 -7 -37 -3
rect -31 -7 -29 -3
rect -14 -7 -12 -3
rect -6 -7 -4 -3
rect 11 -7 13 -3
rect 19 -7 21 -3
rect 40 -7 42 -3
<< ptransistor >>
rect -39 7 -37 11
rect -31 7 -29 11
rect -14 7 -12 11
rect -6 7 -4 11
rect 11 7 13 11
rect 19 7 21 11
rect 40 7 42 11
<< polycontact >>
rect -15 15 -11 19
rect -7 15 -3 19
rect 22 15 26 19
<< ndcontact >>
rect -44 -7 -40 -3
rect -28 -7 -24 -3
rect -19 -7 -15 -3
rect -3 -7 1 -3
rect 6 -7 10 -3
rect 22 -7 26 -3
rect 31 -7 35 -3
rect 47 -7 51 -3
<< pdcontact >>
rect -44 7 -40 11
rect -36 7 -32 11
rect -28 7 -24 11
rect -19 7 -15 11
rect -11 7 -7 11
rect -3 7 1 11
rect 6 7 10 11
rect 14 7 18 11
rect 22 7 26 11
rect 31 7 35 11
rect 47 7 51 11
<< labels >>
rlabel polysilicon -31 13 -29 13 1 SEL
rlabel polysilicon 40 13 42 13 1 SEL
rlabel pdcontact -19 11 -15 11 1 Vdd
rlabel pdcontact -3 11 1 11 1 Vdd
rlabel pdcontact 6 11 10 11 1 Vdd
rlabel pdcontact 22 11 26 11 1 Vdd
rlabel metal1 1 0 1 4 3 Z
rlabel pdcontact -44 11 -40 11 1 Vdd
rlabel pdcontact -28 11 -24 11 1 Vdd
rlabel pdcontact 31 11 35 11 1 Vdd
rlabel metal1 51 -17 51 -14 8 GND
rlabel polysilicon -39 13 -37 13 1 a
rlabel polysilicon 11 13 13 13 1 b
<< end >>
