* SPICE3 file created from nor3.ext - technology: scmos

M1000 a_n2_5# A Vdd w_n10_3# pmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1001 Z C a_6_5# w_n10_3# pmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1002 Z C Gnd Gnd nmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_6_5# B a_n2_5# w_n10_3# pmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1004 Gnd B Z Gnd nmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1005 Z A Gnd Gnd nmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
C0 w_n10_3# B 1.43fF
C1 w_n10_3# A 1.43fF
C2 Z C 0.24fF
C3 Z w_n10_3# 0.38fF
C4 Z B 0.24fF
C5 w_n10_3# C 1.43fF
C6 w_n10_3# Vdd 0.56fF
C7 Gnd Gnd 4.93fF
C8 Z Gnd 4.32fF
C9 Vdd Gnd 4.37fF
C10 C Gnd 2.86fF
C11 B Gnd 2.86fF
C12 A Gnd 2.86fF

VCC    Vdd     GND     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin     A     GND    PWL(   0   0    30N  0    30.1N 2.5   60N  2.5 60.1N  2.5  90N 2.5 90.1N 0 120N 0) 

*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin2     B     GND    PWL(   0   0    30N  0    30.1N 2.5   60N  2.5 60.1N  0  90N 0 90.1N 2.5 120N 2.5)

*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin3     C     GND    PWL(   0   0    30N  0    30.1N 2.5   60N  2.5 60.1N  0  90N 0 90.1N 2.5 120N 2.5) 
 


*     TSTEP TSTOP
*     ----- -----
.TRAN 5N  120N


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
