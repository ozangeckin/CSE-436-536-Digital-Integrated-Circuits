* SPICE3 file created from xor2.ext - technology: scmos

M1000 Z B a_0_n13# Gnd nmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1001 Z B A w_n9_n3# pmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_0_n13# A Gnd Gnd nmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_0_n13# A vdd w_n9_n3# pmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
C0 Z w_n9_n3# 0.75fF
C1 B w_n9_n3# 1.91fF
C2 a_0_n13# w_n9_n3# 1.18fF
C3 A w_n9_n3# 1.91fF
C4 vdd w_n9_n3# 0.56fF
C5 Gnd Gnd 4.65fF
C6 Z Gnd 1.13fF
C7 A Gnd 2.38fF
C8 a_0_n13# Gnd 2.96fF
C9 vdd Gnd 4.09fF
C10 B Gnd 2.38fF

VCC    Vdd     GND     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin     A     GND    PWL(   0   0    30N  0    30.1N 2.5   60N  2.5 60.1N  2.5  90N 2.5 90.1N 2.5 120N 2.5) 

*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin2     B     GND    PWL(   0   2.5    30N  2.5    30.1N 0   60N  0 60.1N  0  90N 0 90.1N 2.5 120N 2.5) 


*     TSTEP TSTOP
*     ----- -----
.TRAN 5N  120N


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END

