magic
tech scmos
timestamp 1639079446
<< nwell >>
rect -9 -3 24 9
<< polysilicon >>
rect -2 5 0 7
rect 15 5 17 7
rect -2 -9 0 1
rect 15 -9 17 1
rect -2 -15 0 -13
rect 15 -15 17 -13
<< ndiffusion >>
rect -3 -13 -2 -9
rect 0 -13 1 -9
rect 14 -13 15 -9
rect 17 -13 18 -9
<< pdiffusion >>
rect -3 1 -2 5
rect 0 1 1 5
rect 14 1 15 5
rect 17 1 18 5
<< metal1 >>
rect -7 9 22 12
rect -7 5 -4 9
rect 1 -2 5 1
rect 1 -6 14 -2
rect 1 -9 5 -6
rect 10 -9 14 -6
rect 18 -9 22 1
rect -7 -17 -4 -13
rect -7 -20 22 -17
<< ntransistor >>
rect -2 -13 0 -9
rect 15 -13 17 -9
<< ptransistor >>
rect -2 1 0 5
rect 15 1 17 5
<< ndcontact >>
rect -7 -13 -3 -9
rect 1 -13 5 -9
rect 10 -13 14 -9
rect 18 -13 22 -9
<< pdcontact >>
rect -7 1 -3 5
rect 1 1 5 5
rect 10 1 14 5
rect 18 1 22 5
<< labels >>
rlabel metal1 22 -6 22 -2 3 Z
rlabel polysilicon 15 7 17 7 1 B
rlabel polysilicon -2 7 0 7 1 A
rlabel pdcontact 10 5 14 5 1 A
rlabel metal1 22 9 22 12 6 vdd
rlabel metal1 22 -20 22 -17 8 Gnd
<< end >>
