* SPICE3 file created from nor2.ext - technology: scmos

M1000 Z A GND Gnd nmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_n11_5# A VDD w_n20_4# pmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1002 GND B Z Gnd nmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1003 Z B a_n11_5# w_n20_4# pmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
C0 w_n20_4# VDD 0.70fF
C1 w_n20_4# Z 0.19fF
C2 w_n20_4# B 1.19fF
C3 Z B 0.24fF
C4 w_n20_4# A 1.19fF
C5 GND Gnd 3.67fF
C6 Z Gnd 2.82fF
C7 VDD Gnd 3.24fF
C8 B Gnd 3.10fF
C9 A Gnd 3.10fF

VCC    Vdd     GND     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin     A     GND    PWL(   0   0    30N  0    30.1N 2.5   60N  2.5 60.1N  2.5  90N 2.5 90.1N 0 120N 0) 

*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin2     B     GND    PWL(   0   0    30N  0    30.1N 2.5   60N  2.5 60.1N  0  90N 0 90.1N 2.5 120N 2.5) 


*     TSTEP TSTOP
*     ----- -----
.TRAN 5N  120N


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
