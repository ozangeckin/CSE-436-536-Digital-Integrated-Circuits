magic
tech scmos
timestamp 1639077816
<< nwell >>
rect -6 1 16 11
<< polysilicon >>
rect 0 8 2 10
rect 8 8 10 10
rect 0 -6 2 4
rect 8 -6 10 4
rect 0 -12 2 -10
rect 8 -12 10 -10
<< ndiffusion >>
rect -1 -10 0 -6
rect 2 -10 8 -6
rect 10 -10 11 -6
<< pdiffusion >>
rect -1 4 0 8
rect 2 4 3 8
rect 7 4 8 8
rect 10 4 11 8
<< metal1 >>
rect -5 12 15 15
rect -5 8 -2 12
rect 12 8 15 12
rect 3 1 7 4
rect 3 -2 15 1
rect 11 -6 15 -2
rect -5 -13 -2 -10
rect -5 -16 15 -13
<< ntransistor >>
rect 0 -10 2 -6
rect 8 -10 10 -6
<< ptransistor >>
rect 0 4 2 8
rect 8 4 10 8
<< ndcontact >>
rect -5 -10 -1 -6
rect 11 -10 15 -6
<< pdcontact >>
rect -5 4 -1 8
rect 3 4 7 8
rect 11 4 15 8
<< labels >>
rlabel metal1 15 -2 15 1 3 Z
rlabel polysilicon 0 10 2 10 1 A
rlabel polysilicon 8 10 10 10 1 B
rlabel metal1 15 12 15 15 6 vdd
rlabel metal1 15 -16 15 -13 8 GND
<< end >>
