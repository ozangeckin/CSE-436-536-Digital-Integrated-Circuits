* SPICE3 file created from nand3.ext - technology: scmos

M1000 a_1_n11# A GND Gnd nmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1001 Z A Vdd w_n8_0# pmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_9_n11# B a_1_n11# Gnd nmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1003 Z C a_9_n11# Gnd nmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1004 Z C Vdd w_n8_0# pmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1005 Vdd B Z w_n8_0# pmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
C0 Z B 0.24fF
C1 B w_n8_0# 1.67fF
C2 A w_n8_0# 1.67fF
C3 Z w_n8_0# 1.13fF
C4 Vdd w_n8_0# 0.85fF
C5 C Z 0.24fF
C6 C w_n8_0# 1.67fF
C7 GND Gnd 4.65fF
C8 Z Gnd 3.57fF
C9 Vdd Gnd 4.37fF
C10 C Gnd 2.62fF
C11 B Gnd 2.62fF
C12 A Gnd 2.62fF

VCC    Vdd     GND     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin     A     GND    PWL(   0   2.5    30N  2.5    30.1N 2.5   60N  2.5 60.1N  2.5  90N 2.5 90.1N 0 120N 0) 

*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin2     B     GND    PWL(   0   0    30N  0    30.1N 2.5   60N  2.5 60.1N  0  90N 0 90.1N 2.5 120N 2.5) 

*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin3     C     GND    PWL(   0   2.5    30N  2.5    30.1N 2.5   60N  2.5 60.1N  0  90N 0 90.1N 2.5 120N 2.5) 


*     TSTEP TSTOP
*     ----- -----
.TRAN 5N  120N


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END

