* SPICE3 file created from /home/ozan/Desktop/integratedCircuit/nand.ext - technology: scmos

M1000 a_n3_n35# A 0 0 nmos w=0.48u l=0.24u
+  ad=0p pd=0u as=0p ps=0u
M1001 F a_n3_n1# 0 0 nmos w=0.48u l=0.24u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_n3_n1# A VDD w_n16_n10# pmos w=0.48u l=0.24u
+  ad=0p pd=0u as=0p ps=0u
M1003 F a_n3_n1# VDD w_n16_n10# pmos w=0.48u l=0.24u
+  ad=0p pd=0u as=0p ps=0u
M1004 VDD B a_n3_n1# w_n16_n10# pmos w=0.48u l=0.24u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_n3_n1# B a_n3_n35# 0 nmos w=0.48u l=0.24u
+  ad=0p pd=0u as=0p ps=0u
C0 B a_n3_n1# 0.13fF
C1 F a_n3_n1# 0.06fF
C2 F 0 0.09fF
C3 VDD F 0.05fF
C4 0 a_n3_n1# 0.05fF
C5 VDD a_n3_n1# 0.07fF
C6 B w_n16_n10# 0.15fF
C7 w_n16_n10# F 0.07fF
C8 w_n16_n10# a_n3_n1# 0.21fF
C9 A B 0.03fF
C10 A a_n3_n1# 0.05fF
C11 w_n16_n10# VDD 0.14fF
C12 A w_n16_n10# 0.15fF
C13 0 0 0.37fF
C14 F 0 0.19fF
C15 VDD 0 0.34fF
C16 a_n3_n1# 0 0.54fF
C17 B 0 0.32fF
C18 A 0 0.32fF
C19 w_n16_n10# 0 0.93fF

* INDEPENDANT VOLTAGE SOURCE
*
*Vname +NODE -NODE VALUE
*----- ----- ----- -----
VCC    VDD     0     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5   
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- --   
VinA     A     0    PWL(   0   0    4N  0    4.1N  2.5   8N  2.5   8.1N  0    12N  0    12.1N  2.5  16N  2.5  16.1N  2.5) 
VinB     B     0    PWL(   0   0    4N  0    4.1N  0     8N  0     8.1N  2.5  12N  2.5  12.1N  2.5  16N  2.5  16.1N  2.5)  

*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  16N


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
