* SPICE3 file created from inverter.ext - technology: scmos

M1000 Z A GND Gnd nmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1001 Z A vdd w_n5_10# pmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
C0 Z w_n5_10# 0.28fF
C1 A w_n5_10# 1.43fF
C2 vdd w_n5_10# 0.56fF
C3 GND Gnd 2.26fF
C4 Z Gnd 1.13fF
C5 vdd Gnd 1.97fF
C6 A Gnd 2.86fF

VCC    Vdd     GND     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin     A     GND    PWL(   0   0    30N  0    30.1N 2.5   60N  2.5 60.1N  2.5  90N 2.5 90.1N 0 120N 0) 


*     TSTEP TSTOP
*     ----- -----
.TRAN 5N  120N


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
