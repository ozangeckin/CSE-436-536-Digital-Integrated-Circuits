magic
tech scmos
timestamp 1639078241
<< nwell >>
rect -20 4 4 14
<< polysilicon >>
rect -13 9 -11 11
rect -5 9 -3 11
rect -13 -5 -11 5
rect -5 -5 -3 5
rect -13 -11 -11 -9
rect -5 -11 -3 -9
<< ndiffusion >>
rect -14 -9 -13 -5
rect -11 -9 -10 -5
rect -6 -9 -5 -5
rect -3 -9 -2 -5
<< pdiffusion >>
rect -14 5 -13 9
rect -11 5 -5 9
rect -3 5 -2 9
<< metal1 >>
rect -18 16 3 19
rect -18 9 -15 16
rect -2 2 2 5
rect -10 -2 2 2
rect -10 -5 -6 -2
rect -18 -12 -15 -9
rect -1 -12 2 -9
rect -18 -15 2 -12
<< ntransistor >>
rect -13 -9 -11 -5
rect -5 -9 -3 -5
<< ptransistor >>
rect -13 5 -11 9
rect -5 5 -3 9
<< ndcontact >>
rect -18 -9 -14 -5
rect -10 -9 -6 -5
rect -2 -9 2 -5
<< pdcontact >>
rect -18 5 -14 9
rect -2 5 2 9
<< labels >>
rlabel polysilicon -13 11 -11 11 1 A
rlabel polysilicon -5 11 -3 11 1 B
rlabel metal1 2 -2 2 2 3 Z
rlabel metal1 3 16 3 19 6 VDD
rlabel metal1 2 -15 2 -12 8 GND
<< end >>
