magic
tech scmos
timestamp 1635249420
<< nwell >>
rect -11 -8 15 13
<< ntransistor >>
rect 0 -22 2 -15
<< ptransistor >>
rect 0 1 2 5
<< ndiffusion >>
rect -1 -22 0 -15
rect 2 -22 3 -15
<< pdiffusion >>
rect -1 1 0 5
rect 2 1 3 5
<< ndcontact >>
rect -5 -22 -1 -15
rect 3 -22 7 -15
<< pdcontact >>
rect -5 1 -1 5
rect 3 1 7 5
<< polysilicon >>
rect 0 5 2 12
rect 0 -15 2 1
rect 0 -25 2 -22
<< polycontact >>
rect -5 -11 0 -5
<< metal1 >>
rect -13 16 17 19
rect -5 5 -2 16
rect -17 -11 -5 -7
rect 4 -7 7 1
rect 4 -10 17 -7
rect 4 -15 7 -10
rect -5 -28 -2 -22
rect -12 -31 14 -28
<< labels >>
rlabel metal1 14 -31 14 -28 8 GND
rlabel metal1 17 16 17 19 6 VDD
rlabel metal1 -17 -11 -17 -7 5 A
rlabel metal1 17 -10 17 -7 5 F
<< end >>
